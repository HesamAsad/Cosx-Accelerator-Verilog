module comp(input[9:0] a,b,output lt);
  assign lt = (a<b);
endmodule
