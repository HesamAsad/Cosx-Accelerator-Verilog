module converter(input[7:0]a,output [9:0]b);
	assign b={2'b00,a};
endmodule
